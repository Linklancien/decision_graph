module main

pub 